module pipeline_wb
(
    input  clk,
          reset
);

  always_ff @ (posedge clk) begin
    
  end
endmodule
